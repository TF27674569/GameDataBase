     