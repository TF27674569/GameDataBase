                           