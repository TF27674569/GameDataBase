                           