!1!3.100~