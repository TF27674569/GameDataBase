       