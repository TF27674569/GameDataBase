                       �          P                            � @   ����������                                                             K   ����    jiaoxue                                                                         